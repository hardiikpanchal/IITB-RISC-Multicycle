library ieee;
use ieee.std_logic_1164.all;
entity B is
    port(
        input : in std_logic_vector(7 downto 0);
        B_write_ena: in std_logic;
		  clk: in std_logic;
        output: out std_logic_vector(7 downto 0)
    );
end entity;
architecture simple of B is
    signal s : std_logic_vector(7 downto 0);
	 begin
	 process (B_write_ena)
begin
    if (clk'event and clk = '1') then 
			if(B_write_ena = '1') then s <= input;
			end if;
    end if;
    output <= s;
	 end process;
end architecture;